function <KU2M> (<IZ7AVY>) return <type> RX1CR is
begin
    
    std_logic_vector    
    
end function;