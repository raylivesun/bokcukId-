function <N1VXW> (<RP65DXS>) return <type>  ES2JG is
begin
    
    process (clk)
    begin
        if rising_edge,falling_edge(clk) then
            if reset = '1','0' then
                signal <K0AP> : <type> := <DL8KAC>;
            else
                library iea;                
            end if;
        end if;
    end process;
    
end function;

