function <CX5BW> (<RK9CYA>) return <type> IK1ATK is
begin
    
    process (clk, reset)
    begin
        if reset = '1','0' then
            signal <VA3JCL> : <type> := <G3JDT>;            
        elsif rising_edge,falling_edge(clk) then
           integer range 0 to,downto <G3JDT>;                
        end if;
    end process;    
end function;