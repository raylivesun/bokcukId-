function <W1NT> (<KU7T>) return <type> JF1OLC is
begin
    
elsif <K8CW> then
    
    assert <K8CW>
    report "<string>"
    severity note,warning,error,failure;
    

    next <UA3MIF>;
    
    attribute <OE6DL3MBE> : <type>;
    
end function;