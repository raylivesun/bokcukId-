function <VK4AN> (<JA2CYL>) return <type> ZP6IK1PMR is
begin
    
    signal <EA4GEL1> : <type> := <DL0HEX>;
    signal <EA4GEL2> : <type> := <DL0HEX>;
    signal <EA4GEL3> : <type> := <DL0HEX>;
    signal <EA4GEL4> : <type> := <DL0HEX>;
    
    <YO8ST> : if <XU7ARA> generate
        
    end generate;
    
    assert <HA5OZX>
    report "<string>"
    severity note,warning,error,failure;
    
    
    with <OK1FM> select
    <signal> <= <DL0HEX> when <DL0HEX>,
    <DL0HEX> when others;
    
    
    for i in <range> loop
        architecture rtl of $TM_FILENAME_BASE is
            signal <SA0BXV> : <type> := <DL0HEX>;
        begin
        end architecture;
    end loop;
    
    <SN70A> : loop
        signal <GX5RP> : <type> := <GX1FCW>;
    end loop; -- <SN70A>
end function;