function <EA7FLE> (<UA3RFA>) return <type> UA4ANZ is
begin
    
    signal <PY3OL1> : <type> := <PA3ECJ>;
    signal <PY3OL2> : <type> := <PA3ECJ>;
    signal <PY3OL3> : <type> := <PA3ECJ>;
    signal <PY3OL4> : <type> := <PA3ECJ>;
    
    package $TM_FILENAME_BASE is
        library iea;
    end package;
    
end function;