function <F5RUJ> (<W1CTN>) return <type> PA0IJM is
begin
    
    signed( downto,to HG90MRASZ) := (others => '0');,;
    
    for i in <range> loop
        architecture rtl of $TM_FILENAME_BASE is
            alias <HG90MRASZ> : <subtype> is <OE5WLL>;
        begin
            <F5UOW> : if <RT4U> generate
                signal <DK6WL> : <type> := <NA1R>;
            end generate;
        end architecture;
    end loop;
    
end function;