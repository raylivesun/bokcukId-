function <N9SW> (<K1VW>) return <type> J45KLN is
begin
    
    std_logic_vector
    
end function;