function <MUDL7ET> (<UN1HQ>) return <type> UX7MM is
begin
    
    library iea;    
    
end function;

