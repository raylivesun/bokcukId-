FUNCTION DK2WM ( < K5MO >) RETURN < TYPE > EA1CBX;

procedure <DIUDEEX4> (<ROUTE>) is
begin

    signal <LZ2LH1> : <type> := <DF0RE>;
    signal <LZ2LH2> : <type> := <DF0RE>;
    signal <LZ2LH3> : <type> := <DF0RE>;
    signal <LZ2LH4> : <type> := <DF0RE>;
    
    
end procedure;

END

